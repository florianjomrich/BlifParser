`timescale 1ns / 1ps 
 
module TEST; 
 
// Inputs 
reg \A2.PAD.PAD ;
reg \A1.PAD.PAD ;
reg \A3.PAD.PAD ;
reg \A0.PAD.PAD ;
reg \B3.PAD.PAD ;
reg \B2.PAD.PAD ;
reg \my_clk.PAD.PAD ;
reg \CIN.PAD.PAD ;
reg \B0.PAD.PAD ;
reg \B1.PAD.PAD ;

// Outputs 
wire \S2_FINAL_OUTPUT.OUTBUF.OUT ;
wire \S0_FINAL_OUTPUT.OUTBUF.OUT ;
wire \S1_FINAL_OUTPUT.OUTBUF.OUT ;
wire \S3_FINAL_OUTPUT.OUTBUF.OUT ;
wire \COUT_FINAL_OUTPUT.OUTBUF.OUT ;
wire [4:0] sum;
 
// Instantiate the Unit Under Test (UUT) 
 
helloWorld uut (
.\A2.PAD.PAD (\A2.PAD.PAD ),
.\A1.PAD.PAD (\A1.PAD.PAD ),
.\A3.PAD.PAD (\A3.PAD.PAD ),
.\A0.PAD.PAD (\A0.PAD.PAD ),
.\B3.PAD.PAD (\B3.PAD.PAD ),
.\B2.PAD.PAD (\B2.PAD.PAD ),
.\my_clk.PAD.PAD (\my_clk.PAD.PAD ),
.\CIN.PAD.PAD (\CIN.PAD.PAD ),
.\B0.PAD.PAD (\B0.PAD.PAD ),
.\B1.PAD.PAD (\B1.PAD.PAD ),
.\S2_FINAL_OUTPUT.OUTBUF.OUT (\S2_FINAL_OUTPUT.OUTBUF.OUT ),
.\S0_FINAL_OUTPUT.OUTBUF.OUT (\S0_FINAL_OUTPUT.OUTBUF.OUT ),
.\S1_FINAL_OUTPUT.OUTBUF.OUT (\S1_FINAL_OUTPUT.OUTBUF.OUT ),
.\S3_FINAL_OUTPUT.OUTBUF.OUT (\S3_FINAL_OUTPUT.OUTBUF.OUT ),
.\COUT_FINAL_OUTPUT.OUTBUF.OUT (\COUT_FINAL_OUTPUT.OUTBUF.OUT )
);

initial begin
// Initialize Inputs
\A2.PAD.PAD  = 0;
\A1.PAD.PAD  = 0;
\A3.PAD.PAD  = 0;
\A0.PAD.PAD  = 0;
\B3.PAD.PAD  = 0;
\B2.PAD.PAD  = 0;
\my_clk.PAD.PAD  = 0;
\CIN.PAD.PAD  = 0;
\B0.PAD.PAD  = 0;
\B1.PAD.PAD  = 0;


// Wait 100 ns for global reset to finish
	#100;

	// Add stimulus here
	\A0.PAD.PAD =1;
	#100;
	\B0.PAD.PAD  = 1;
	\B1.PAD.PAD  = 1;
	#100;
	\A3.PAD.PAD =1;
	\B2.PAD.PAD =1;

end

assign sum = {\COUT_FINAL_OUTPUT.OUTBUF.OUT ,\S3_FINAL_OUTPUT.OUTBUF.OUT ,\S2_FINAL_OUTPUT.OUTBUF.OUT , \S1_FINAL_OUTPUT.OUTBUF.OUT ,\S0_FINAL_OUTPUT.OUTBUF.OUT };


endmodule