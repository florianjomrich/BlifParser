//    Xilinx Proprietary Primitive Cell X_ONE for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verplex_libs/data/simprims/X_ONE.v,v 1.4.198.3 2004/09/28 20:47:46 wloo Exp $
//

`celldefine
`timescale 1 ps/1 ps

module X_ONE (O);

  output O;

  assign O = 1'b1;

endmodule
