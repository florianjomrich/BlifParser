// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verplex_libs/data/simprims/X_PPC405.v,v 1.7.144.3 2004/09/28 20:47:46 wloo Exp $

/*

		: Power PC

*/

`timescale  1 ps / 1 ps

module X_PPC405 (
		C405CPMCORESLEEPREQ,
		C405CPMMSRCE,
		C405CPMMSREE,
		C405CPMTIMERIRQ,
		C405CPMTIMERRESETREQ,
		C405DBGMSRWE,
		C405DBGSTOPACK,
		C405DBGWBCOMPLETE,
		C405DBGWBFULL,
		C405DBGWBIAR,
		C405DCRABUS,
		C405DCRDBUSOUT,
		C405DCRREAD,
		C405DCRWRITE,
		C405JTGCAPTUREDR,
		C405JTGEXTEST,
		C405JTGPGMOUT,
		C405JTGSHIFTDR,
		C405JTGTDO,
		C405JTGTDOEN,
		C405JTGUPDATEDR,
		C405PLBDCUABORT,
		C405PLBDCUABUS,
		C405PLBDCUBE,
		C405PLBDCUCACHEABLE,
		C405PLBDCUGUARDED,
		C405PLBDCUPRIORITY,
		C405PLBDCUREQUEST,
		C405PLBDCURNW,
		C405PLBDCUSIZE2,
		C405PLBDCUU0ATTR,
		C405PLBDCUWRDBUS,
		C405PLBDCUWRITETHRU,
		C405PLBICUABORT,
		C405PLBICUABUS,
		C405PLBICUCACHEABLE,
		C405PLBICUPRIORITY,
		C405PLBICUREQUEST,
		C405PLBICUSIZE,
		C405PLBICUU0ATTR,
		C405RSTCHIPRESETREQ,
		C405RSTCORERESETREQ,
		C405RSTSYSRESETREQ,
		C405TRCCYCLE,
		C405TRCEVENEXECUTIONSTATUS,
		C405TRCODDEXECUTIONSTATUS,
		C405TRCTRACESTATUS,
		C405TRCTRIGGEREVENTOUT,
		C405TRCTRIGGEREVENTTYPE,
		C405XXXMACHINECHECK,
		DSOCMBRAMABUS,
		DSOCMBRAMBYTEWRITE,
		DSOCMBRAMEN,
		DSOCMBRAMWRDBUS,
		DSOCMBUSY,
		ISOCMBRAMEN,
		ISOCMBRAMEVENWRITEEN,
		ISOCMBRAMODDWRITEEN,
		ISOCMBRAMRDABUS,
		ISOCMBRAMWRABUS,
		ISOCMBRAMWRDBUS,

		BRAMDSOCMCLK,
		BRAMDSOCMRDDBUS,
		BRAMISOCMCLK,
		BRAMISOCMRDDBUS,
		CPMC405CLOCK,
		CPMC405CORECLKINACTIVE,
		CPMC405CPUCLKEN,
		CPMC405JTAGCLKEN,
		CPMC405TIMERCLKEN,
		CPMC405TIMERTICK,
		DBGC405DEBUGHALT,
		DBGC405EXTBUSHOLDACK,
		DBGC405UNCONDDEBUGEVENT,
		DCRC405ACK,
		DCRC405DBUSIN,
		DSARCVALUE,
		DSCNTLVALUE,
		EICC405CRITINPUTIRQ,
		EICC405EXTINPUTIRQ,
		ISARCVALUE,
		ISCNTLVALUE,
		JTGC405BNDSCANTDO,
		JTGC405TCK,
		JTGC405TDI,
		JTGC405TMS,
		JTGC405TRSTNEG,
		MCBCPUCLKEN,
		MCBJTAGEN,
		MCBTIMEREN,
		MCPPCRST,
		PLBC405DCUADDRACK,
		PLBC405DCUBUSY,
		PLBC405DCUERR,
		PLBC405DCURDDACK,
		PLBC405DCURDDBUS,
		PLBC405DCURDWDADDR,
		PLBC405DCUSSIZE1,
		PLBC405DCUWRDACK,
		PLBC405ICUADDRACK,
		PLBC405ICUBUSY,
		PLBC405ICUERR,
		PLBC405ICURDDACK,
		PLBC405ICURDDBUS,
		PLBC405ICURDWDADDR,
		PLBC405ICUSSIZE1,
		PLBCLK,
		RSTC405RESETCHIP,
		RSTC405RESETCORE,
		RSTC405RESETSYS,
		TIEC405DETERMINISTICMULT,
		TIEC405DISOPERANDFWD,
		TIEC405MMUEN,
		TIEDSOCMDCRADDR,
		TIEISOCMDCRADDR,
		TRCC405TRACEDISABLE,
		TRCC405TRIGGEREVENTIN
);

parameter in_delay=0;
parameter out_delay=0;
parameter PPCUSER = 4'b0000;

output		C405CPMCORESLEEPREQ;
output		C405CPMMSRCE;
output		C405CPMMSREE;
output		C405CPMTIMERIRQ;
output		C405CPMTIMERRESETREQ;
output		C405DBGMSRWE;
output		C405DBGSTOPACK;
output		C405DBGWBCOMPLETE;
output		C405DBGWBFULL;
output	[0:29]	C405DBGWBIAR;
output	[0:9]	C405DCRABUS;
output	[0:31]	C405DCRDBUSOUT;
output		C405DCRREAD;
output		C405DCRWRITE;
output		C405JTGCAPTUREDR;
output		C405JTGEXTEST;
output		C405JTGPGMOUT;
output		C405JTGSHIFTDR;
output		C405JTGTDO;
output		C405JTGTDOEN;
output		C405JTGUPDATEDR;
output		C405PLBDCUABORT;
output	[0:31]	C405PLBDCUABUS;
output	[0:7]	C405PLBDCUBE;
output		C405PLBDCUCACHEABLE;
output		C405PLBDCUGUARDED;
output	[0:1]	C405PLBDCUPRIORITY;
output		C405PLBDCUREQUEST;
output		C405PLBDCURNW;
output		C405PLBDCUSIZE2;
output		C405PLBDCUU0ATTR;
output	[0:63]	C405PLBDCUWRDBUS;
output		C405PLBDCUWRITETHRU;
output		C405PLBICUABORT;
output	[0:29]	C405PLBICUABUS;
output		C405PLBICUCACHEABLE;
output	[0:1]	C405PLBICUPRIORITY;
output		C405PLBICUREQUEST;
output	[2:3]	C405PLBICUSIZE;
output		C405PLBICUU0ATTR;
output		C405RSTCHIPRESETREQ;
output		C405RSTCORERESETREQ;
output		C405RSTSYSRESETREQ;
output		C405TRCCYCLE;
output	[0:1]	C405TRCEVENEXECUTIONSTATUS;
output	[0:1]	C405TRCODDEXECUTIONSTATUS;
output	[0:3]	C405TRCTRACESTATUS;
output		C405TRCTRIGGEREVENTOUT;
output	[0:10]	C405TRCTRIGGEREVENTTYPE;
output		C405XXXMACHINECHECK;
output	[8:29]	DSOCMBRAMABUS;
output	[0:3]	DSOCMBRAMBYTEWRITE;
output		DSOCMBRAMEN;
output	[0:31]	DSOCMBRAMWRDBUS;
output		DSOCMBUSY;
output		ISOCMBRAMEN;
output		ISOCMBRAMEVENWRITEEN;
output		ISOCMBRAMODDWRITEEN;
output	[8:28]	ISOCMBRAMRDABUS;
output	[8:28]	ISOCMBRAMWRABUS;
output	[0:31]	ISOCMBRAMWRDBUS;

input		BRAMDSOCMCLK;
input	[0:31]	BRAMDSOCMRDDBUS;
input		BRAMISOCMCLK;
input	[0:63]	BRAMISOCMRDDBUS;
input		CPMC405CLOCK;
input		CPMC405CORECLKINACTIVE;
input		CPMC405CPUCLKEN;
input		CPMC405JTAGCLKEN;
input		CPMC405TIMERCLKEN;
input		CPMC405TIMERTICK;
input		DBGC405DEBUGHALT;
input		DBGC405EXTBUSHOLDACK;
input		DBGC405UNCONDDEBUGEVENT;
input		DCRC405ACK;
input	[0:31]	DCRC405DBUSIN;
input	[0:7]	DSARCVALUE;
input	[0:7]	DSCNTLVALUE;
input		EICC405CRITINPUTIRQ;
input		EICC405EXTINPUTIRQ;
input	[0:7]	ISARCVALUE;
input	[0:7]	ISCNTLVALUE;
input		JTGC405BNDSCANTDO;
input		JTGC405TCK;
input		JTGC405TDI;
input		JTGC405TMS;
input		JTGC405TRSTNEG;
input		MCBCPUCLKEN;
input		MCBJTAGEN;
input		MCBTIMEREN;
input		MCPPCRST;
input		PLBC405DCUADDRACK;
input		PLBC405DCUBUSY;
input		PLBC405DCUERR;
input		PLBC405DCURDDACK;
input	[0:63]	PLBC405DCURDDBUS;
input	[1:3]	PLBC405DCURDWDADDR;
input		PLBC405DCUSSIZE1;
input		PLBC405DCUWRDACK;
input		PLBC405ICUADDRACK;
input		PLBC405ICUBUSY;
input		PLBC405ICUERR;
input		PLBC405ICURDDACK;
input	[0:63]	PLBC405ICURDDBUS;
input	[1:3]	PLBC405ICURDWDADDR;
input		PLBC405ICUSSIZE1;
input		PLBCLK;
input		RSTC405RESETCHIP;
input		RSTC405RESETCORE;
input		RSTC405RESETSYS;
input		TIEC405DETERMINISTICMULT;
input		TIEC405DISOPERANDFWD;
input		TIEC405MMUEN;
input	[0:7]	TIEDSOCMDCRADDR;
input	[0:7]	TIEISOCMDCRADDR;
input		TRCC405TRACEDISABLE;
input		TRCC405TRIGGEREVENTIN;
   
endmodule
