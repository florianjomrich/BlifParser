//    Xilinx Proprietary Primitive Cell X_MUXDDR for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verplex_libs/data/simprims/X_MUXDDR.v,v 1.4.198.3 2004/09/28 20:47:46 wloo Exp $
//

`celldefine
`timescale 1 ps/1 ps


module X_MUXDDR (O, CE, CLK0, CLK1, I0, I1);

    output O;

    input  CE, CLK0, CLK1, I0, I1;

endmodule
