`timescale 1ns / 1ps 
 
module TEST; 
 
// Inputs 
reg \key<173>.PAD.PAD ;
reg \key<89>.PAD.PAD ;
reg \key<8>.PAD.PAD ;
reg \key<183>.PAD.PAD ;
reg \key<108>.PAD.PAD ;
reg \key<99>.PAD.PAD ;
reg \key<174>.PAD.PAD ;
reg \key<9>.PAD.PAD ;
reg \key<184>.PAD.PAD ;
reg \key<107>.PAD.PAD ;
reg \key<39>.PAD.PAD ;
reg \key<19>.PAD.PAD ;
reg \key<77>.PAD.PAD ;
reg \key<185>.PAD.PAD ;
reg \key<97>.PAD.PAD ;
reg \key<199>.PAD.PAD ;
reg \key<171>.PAD.PAD ;
reg \key<59>.PAD.PAD ;
reg \key<38>.PAD.PAD ;
reg \key<172>.PAD.PAD ;
reg \key<18>.PAD.PAD ;
reg \key<78>.PAD.PAD ;
reg \key<186>.PAD.PAD ;
reg \key<109>.PAD.PAD ;
reg \key<98>.PAD.PAD ;
reg \key<79>.PAD.PAD ;
reg \key<119>.PAD.PAD ;
reg \key<58>.PAD.PAD ;
reg \key<187>.PAD.PAD ;
reg \key<47>.PAD.PAD ;
reg \key<75>.PAD.PAD ;
reg \key<4>.PAD.PAD ;
reg \key<37>.PAD.PAD ;
reg \key<177>.PAD.PAD ;
reg \key<85>.PAD.PAD ;
reg \key<118>.PAD.PAD ;
reg \key<197>.PAD.PAD ;
reg \key<104>.PAD.PAD ;
reg \key<188>.PAD.PAD ;
reg \key<5>.PAD.PAD ;
reg \key<76>.PAD.PAD ;
reg \key<46>.PAD.PAD ;
reg \key<36>.PAD.PAD ;
reg \key<86>.PAD.PAD ;
reg \key<178>.PAD.PAD ;
reg \key<117>.PAD.PAD ;
reg \key<198>.PAD.PAD ;
reg \key<45>.PAD.PAD ;
reg \key<103>.PAD.PAD ;
reg \key<6>.PAD.PAD ;
reg \key<49>.PAD.PAD ;
reg \key<211>.PAD.PAD ;
reg \key<73>.PAD.PAD ;
reg \key<189>.PAD.PAD ;
reg \key<87>.PAD.PAD ;
reg \key<35>.PAD.PAD ;
reg \key<175>.PAD.PAD ;
reg \key<116>.PAD.PAD ;
reg \key<34>.PAD.PAD ;
reg \key<195>.PAD.PAD ;
reg \key<106>.PAD.PAD ;
reg \key<48>.PAD.PAD ;
reg \key<7>.PAD.PAD ;
reg \key<210>.PAD.PAD ;
reg \key<74>.PAD.PAD ;
reg \key<176>.PAD.PAD ;
reg \key<88>.PAD.PAD ;
reg \key<33>.PAD.PAD ;
reg \key<115>.PAD.PAD ;
reg \key<196>.PAD.PAD ;
reg \key<105>.PAD.PAD ;
reg \key<213>.PAD.PAD ;
reg \key<42>.PAD.PAD ;
reg \key<127>.PAD.PAD ;
reg \key<32>.PAD.PAD ;
reg \key<227>.PAD.PAD ;
reg \key<0>.PAD.PAD ;
reg \key<52>.PAD.PAD ;
reg \key<62>.PAD.PAD ;
reg \key<41>.PAD.PAD ;
reg \key<128>.PAD.PAD ;
reg \key<226>.PAD.PAD ;
reg \key<31>.PAD.PAD ;
reg \key<212>.PAD.PAD ;
reg \key<1>.PAD.PAD ;
reg \key<51>.PAD.PAD ;
reg \key<61>.PAD.PAD ;
reg \key<139>.PAD.PAD ;
reg \key<44>.PAD.PAD ;
reg \key<215>.PAD.PAD ;
reg \key<225>.PAD.PAD ;
reg \key<129>.PAD.PAD ;
reg \key<30>.PAD.PAD ;
reg \key<179>.PAD.PAD ;
reg \key<2>.PAD.PAD ;
reg \key<50>.PAD.PAD ;
reg \global_reset.PAD.PAD ;
reg \key<64>.PAD.PAD ;
reg \key<43>.PAD.PAD ;
reg \key<214>.PAD.PAD ;
reg \key<224>.PAD.PAD ;
reg \encrypt<0>.PAD.PAD ;
reg \key<3>.PAD.PAD ;
reg \key<63>.PAD.PAD ;
reg \key<57>.PAD.PAD ;
reg \count<0>.PAD.PAD ;
reg \key<217>.PAD.PAD ;
reg \key<66>.PAD.PAD ;
reg \key<237>.PAD.PAD ;
reg \key<56>.PAD.PAD ;
reg \count<1>.PAD.PAD ;
reg \key<216>.PAD.PAD ;
reg \key<65>.PAD.PAD ;
reg \key<236>.PAD.PAD ;
reg \key<55>.PAD.PAD ;
reg \key<229>.PAD.PAD ;
reg \key<40>.PAD.PAD ;
reg \key<69>.PAD.PAD ;
reg \key<219>.PAD.PAD ;
reg \key<239>.PAD.PAD ;
reg \key<54>.PAD.PAD ;
reg \key<249>.PAD.PAD ;
reg \start<0>.PAD.PAD ;
reg \my_clk.PAD.PAD ;
reg \key<228>.PAD.PAD ;
reg \key<68>.PAD.PAD ;
reg \key<218>.PAD.PAD ;
reg \key<238>.PAD.PAD ;
reg \key<67>.PAD.PAD ;
reg \key<248>.PAD.PAD ;
reg \key<53>.PAD.PAD ;
reg \key<208>.PAD.PAD ;
reg \key<244>.PAD.PAD ;
reg \key<132>.PAD.PAD ;
reg \key<230>.PAD.PAD ;
reg \key<146>.PAD.PAD ;
reg \key<245>.PAD.PAD ;
reg \key<209>.PAD.PAD ;
reg \key<159>.PAD.PAD ;
reg \key<131>.PAD.PAD ;
reg \key<231>.PAD.PAD ;
reg \key<145>.PAD.PAD ;
reg \key<246>.PAD.PAD ;
reg \key<134>.PAD.PAD ;
reg \key<144>.PAD.PAD ;
reg \key<247>.PAD.PAD ;
reg \key<133>.PAD.PAD ;
reg \key<143>.PAD.PAD ;
reg \key<156>.PAD.PAD ;
reg \key<254>.PAD.PAD ;
reg \count<3>.PAD.PAD ;
reg \key<240>.PAD.PAD ;
reg \key<220>.PAD.PAD ;
reg \key<136>.PAD.PAD ;
reg \key<234>.PAD.PAD ;
reg \key<155>.PAD.PAD ;
reg \key<169>.PAD.PAD ;
reg \key<255>.PAD.PAD ;
reg \count<2>.PAD.PAD ;
reg \key<241>.PAD.PAD ;
reg \key<221>.PAD.PAD ;
reg \key<235>.PAD.PAD ;
reg \key<20>.PAD.PAD ;
reg \key<149>.PAD.PAD ;
reg \key<135>.PAD.PAD ;
reg \key<252>.PAD.PAD ;
reg \key<168>.PAD.PAD ;
reg \key<158>.PAD.PAD ;
reg \key<242>.PAD.PAD ;
reg \key<138>.PAD.PAD ;
reg \key<222>.PAD.PAD ;
reg \key<232>.PAD.PAD ;
reg \key<148>.PAD.PAD ;
reg \key<253>.PAD.PAD ;
reg \key<60>.PAD.PAD ;
reg \key<157>.PAD.PAD ;
reg \key<167>.PAD.PAD ;
reg \key<243>.PAD.PAD ;
reg \key<137>.PAD.PAD ;
reg \key<223>.PAD.PAD ;
reg \key<233>.PAD.PAD ;
reg \key<147>.PAD.PAD ;
reg \key<111>.PAD.PAD ;
reg \key<125>.PAD.PAD ;
reg \key<92>.PAD.PAD ;
reg \key<194>.PAD.PAD ;
reg \key<23>.PAD.PAD ;
reg \key<24>.PAD.PAD ;
reg \key<82>.PAD.PAD ;
reg \key<166>.PAD.PAD ;
reg \key<250>.PAD.PAD ;
reg \key<200>.PAD.PAD ;
reg \key<72>.PAD.PAD ;
reg \key<152>.PAD.PAD ;
reg \key<10>.PAD.PAD ;
reg \key<112>.PAD.PAD ;
reg \key<91>.PAD.PAD ;
reg \key<126>.PAD.PAD ;
reg \key<193>.PAD.PAD ;
reg \key<25>.PAD.PAD ;
reg \key<165>.PAD.PAD ;
reg \key<201>.PAD.PAD ;
reg \key<251>.PAD.PAD ;
reg \key<81>.PAD.PAD ;
reg \key<71>.PAD.PAD ;
reg \key<151>.PAD.PAD ;
reg \key<123>.PAD.PAD ;
reg \key<11>.PAD.PAD ;
reg \key<21>.PAD.PAD ;
reg \key<90>.PAD.PAD ;
reg \key<113>.PAD.PAD ;
reg \key<202>.PAD.PAD ;
reg \key<192>.PAD.PAD ;
reg \key<84>.PAD.PAD ;
reg \key<164>.PAD.PAD ;
reg \key<70>.PAD.PAD ;
reg \key<154>.PAD.PAD ;
reg \key<124>.PAD.PAD ;
reg \key<114>.PAD.PAD ;
reg \key<12>.PAD.PAD ;
reg \key<22>.PAD.PAD ;
reg \key<203>.PAD.PAD ;
reg \key<163>.PAD.PAD ;
reg \key<191>.PAD.PAD ;
reg \key<83>.PAD.PAD ;
reg \key<153>.PAD.PAD ;
reg \key<13>.PAD.PAD ;
reg \key<170>.PAD.PAD ;
reg \key<142>.PAD.PAD ;
reg \key<121>.PAD.PAD ;
reg \key<180>.PAD.PAD ;
reg \key<96>.PAD.PAD ;
reg \key<14>.PAD.PAD ;
reg \key<101>.PAD.PAD ;
reg \key<162>.PAD.PAD ;
reg \key<190>.PAD.PAD ;
reg \key<28>.PAD.PAD ;
reg \key<204>.PAD.PAD ;
reg \key<141>.PAD.PAD ;
reg \key<95>.PAD.PAD ;
reg \key<122>.PAD.PAD ;
reg \key<102>.PAD.PAD ;
reg \key<15>.PAD.PAD ;
reg \key<161>.PAD.PAD ;
reg \key<205>.PAD.PAD ;
reg \key<29>.PAD.PAD ;
reg \key<160>.PAD.PAD ;
reg \key<140>.PAD.PAD ;
reg \key<94>.PAD.PAD ;
reg \key<130>.PAD.PAD ;
reg \key<182>.PAD.PAD ;
reg \key<150>.PAD.PAD ;
reg \key<16>.PAD.PAD ;
reg \key<80>.PAD.PAD ;
reg \key<206>.PAD.PAD ;
reg \key<26>.PAD.PAD ;
reg \key<110>.PAD.PAD ;
reg \key<181>.PAD.PAD ;
reg \key<93>.PAD.PAD ;
reg \key<120>.PAD.PAD ;
reg \key<100>.PAD.PAD ;
reg \key<17>.PAD.PAD ;
reg \key<27>.PAD.PAD ;
reg \key<207>.PAD.PAD ;

// Outputs 
wire \KSi<19>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<163>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<17>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<55>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<37>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<26>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<136>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<174>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<67>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<6>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<77>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<15>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<108>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<13>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<86>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<150>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<85>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<157>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<113>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<41>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<110>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<104>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<83>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<89>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<11>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<7>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<164>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<179>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<109>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<173>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<155>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<31>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<123>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<44>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<84>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \new_count<2>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<5>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<118>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<141>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<165>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<130>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<162>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<33>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<161>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<154>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<64>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<78>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<170>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<1>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<135>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<95>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<139>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<49>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<12>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<146>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<61>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \data_ready<0>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<34>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<62>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<24>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<53>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<0>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<125>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<22>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<9>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<48>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<111>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<70>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<74>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<79>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<58>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<2>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<29>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<148>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<186>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<68>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<99>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<190>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<105>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<119>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<35>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<133>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<188>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<158>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<115>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<46>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<93>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<73>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<28>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<143>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<54>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<18>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<177>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<106>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<98>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<30>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<142>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<167>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<3>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<60>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<181>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<39>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \new_count<0>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<132>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<16>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<191>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<45>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<116>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<47>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<81>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<100>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<168>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<59>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<121>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<72>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<159>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<14>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<25>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<82>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<90>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<36>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<97>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<175>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<134>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<151>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<10>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<80>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<138>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<169>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<149>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<176>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<140>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<71>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<153>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<145>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<124>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<8>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<172>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<40>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<96>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<75>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<103>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<122>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<129>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<183>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<156>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<4>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<38>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<128>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<107>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<23>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<88>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<185>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<57>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<187>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<50>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<160>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<144>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<32>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<21>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<102>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<137>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<131>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \new_count<1>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<152>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<94>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<182>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<189>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<56>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<52>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<171>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<87>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<51>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<65>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<114>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<76>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<126>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<91>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<92>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<117>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<27>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<66>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<69>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<101>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<178>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<43>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<112>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<166>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<180>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<127>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<147>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<184>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<20>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<42>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \new_count<3>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<120>_FINAL_OUTPUT.OUTBUF.OUT ;
wire \KSi<63>_FINAL_OUTPUT.OUTBUF.OUT ;
 
// Instantiate the Unit Under Test (UUT) 
 
HelloWorld uut (
.\key<173>.PAD.PAD (\key<173>.PAD.PAD ),
.\key<89>.PAD.PAD (\key<89>.PAD.PAD ),
.\key<8>.PAD.PAD (\key<8>.PAD.PAD ),
.\key<183>.PAD.PAD (\key<183>.PAD.PAD ),
.\key<108>.PAD.PAD (\key<108>.PAD.PAD ),
.\key<99>.PAD.PAD (\key<99>.PAD.PAD ),
.\key<174>.PAD.PAD (\key<174>.PAD.PAD ),
.\key<9>.PAD.PAD (\key<9>.PAD.PAD ),
.\key<184>.PAD.PAD (\key<184>.PAD.PAD ),
.\key<107>.PAD.PAD (\key<107>.PAD.PAD ),
.\key<39>.PAD.PAD (\key<39>.PAD.PAD ),
.\key<19>.PAD.PAD (\key<19>.PAD.PAD ),
.\key<77>.PAD.PAD (\key<77>.PAD.PAD ),
.\key<185>.PAD.PAD (\key<185>.PAD.PAD ),
.\key<97>.PAD.PAD (\key<97>.PAD.PAD ),
.\key<199>.PAD.PAD (\key<199>.PAD.PAD ),
.\key<171>.PAD.PAD (\key<171>.PAD.PAD ),
.\key<59>.PAD.PAD (\key<59>.PAD.PAD ),
.\key<38>.PAD.PAD (\key<38>.PAD.PAD ),
.\key<172>.PAD.PAD (\key<172>.PAD.PAD ),
.\key<18>.PAD.PAD (\key<18>.PAD.PAD ),
.\key<78>.PAD.PAD (\key<78>.PAD.PAD ),
.\key<186>.PAD.PAD (\key<186>.PAD.PAD ),
.\key<109>.PAD.PAD (\key<109>.PAD.PAD ),
.\key<98>.PAD.PAD (\key<98>.PAD.PAD ),
.\key<79>.PAD.PAD (\key<79>.PAD.PAD ),
.\key<119>.PAD.PAD (\key<119>.PAD.PAD ),
.\key<58>.PAD.PAD (\key<58>.PAD.PAD ),
.\key<187>.PAD.PAD (\key<187>.PAD.PAD ),
.\key<47>.PAD.PAD (\key<47>.PAD.PAD ),
.\key<75>.PAD.PAD (\key<75>.PAD.PAD ),
.\key<4>.PAD.PAD (\key<4>.PAD.PAD ),
.\key<37>.PAD.PAD (\key<37>.PAD.PAD ),
.\key<177>.PAD.PAD (\key<177>.PAD.PAD ),
.\key<85>.PAD.PAD (\key<85>.PAD.PAD ),
.\key<118>.PAD.PAD (\key<118>.PAD.PAD ),
.\key<197>.PAD.PAD (\key<197>.PAD.PAD ),
.\key<104>.PAD.PAD (\key<104>.PAD.PAD ),
.\key<188>.PAD.PAD (\key<188>.PAD.PAD ),
.\key<5>.PAD.PAD (\key<5>.PAD.PAD ),
.\key<76>.PAD.PAD (\key<76>.PAD.PAD ),
.\key<46>.PAD.PAD (\key<46>.PAD.PAD ),
.\key<36>.PAD.PAD (\key<36>.PAD.PAD ),
.\key<86>.PAD.PAD (\key<86>.PAD.PAD ),
.\key<178>.PAD.PAD (\key<178>.PAD.PAD ),
.\key<117>.PAD.PAD (\key<117>.PAD.PAD ),
.\key<198>.PAD.PAD (\key<198>.PAD.PAD ),
.\key<45>.PAD.PAD (\key<45>.PAD.PAD ),
.\key<103>.PAD.PAD (\key<103>.PAD.PAD ),
.\key<6>.PAD.PAD (\key<6>.PAD.PAD ),
.\key<49>.PAD.PAD (\key<49>.PAD.PAD ),
.\key<211>.PAD.PAD (\key<211>.PAD.PAD ),
.\key<73>.PAD.PAD (\key<73>.PAD.PAD ),
.\key<189>.PAD.PAD (\key<189>.PAD.PAD ),
.\key<87>.PAD.PAD (\key<87>.PAD.PAD ),
.\key<35>.PAD.PAD (\key<35>.PAD.PAD ),
.\key<175>.PAD.PAD (\key<175>.PAD.PAD ),
.\key<116>.PAD.PAD (\key<116>.PAD.PAD ),
.\key<34>.PAD.PAD (\key<34>.PAD.PAD ),
.\key<195>.PAD.PAD (\key<195>.PAD.PAD ),
.\key<106>.PAD.PAD (\key<106>.PAD.PAD ),
.\key<48>.PAD.PAD (\key<48>.PAD.PAD ),
.\key<7>.PAD.PAD (\key<7>.PAD.PAD ),
.\key<210>.PAD.PAD (\key<210>.PAD.PAD ),
.\key<74>.PAD.PAD (\key<74>.PAD.PAD ),
.\key<176>.PAD.PAD (\key<176>.PAD.PAD ),
.\key<88>.PAD.PAD (\key<88>.PAD.PAD ),
.\key<33>.PAD.PAD (\key<33>.PAD.PAD ),
.\key<115>.PAD.PAD (\key<115>.PAD.PAD ),
.\key<196>.PAD.PAD (\key<196>.PAD.PAD ),
.\key<105>.PAD.PAD (\key<105>.PAD.PAD ),
.\key<213>.PAD.PAD (\key<213>.PAD.PAD ),
.\key<42>.PAD.PAD (\key<42>.PAD.PAD ),
.\key<127>.PAD.PAD (\key<127>.PAD.PAD ),
.\key<32>.PAD.PAD (\key<32>.PAD.PAD ),
.\key<227>.PAD.PAD (\key<227>.PAD.PAD ),
.\key<0>.PAD.PAD (\key<0>.PAD.PAD ),
.\key<52>.PAD.PAD (\key<52>.PAD.PAD ),
.\key<62>.PAD.PAD (\key<62>.PAD.PAD ),
.\key<41>.PAD.PAD (\key<41>.PAD.PAD ),
.\key<128>.PAD.PAD (\key<128>.PAD.PAD ),
.\key<226>.PAD.PAD (\key<226>.PAD.PAD ),
.\key<31>.PAD.PAD (\key<31>.PAD.PAD ),
.\key<212>.PAD.PAD (\key<212>.PAD.PAD ),
.\key<1>.PAD.PAD (\key<1>.PAD.PAD ),
.\key<51>.PAD.PAD (\key<51>.PAD.PAD ),
.\key<61>.PAD.PAD (\key<61>.PAD.PAD ),
.\key<139>.PAD.PAD (\key<139>.PAD.PAD ),
.\key<44>.PAD.PAD (\key<44>.PAD.PAD ),
.\key<215>.PAD.PAD (\key<215>.PAD.PAD ),
.\key<225>.PAD.PAD (\key<225>.PAD.PAD ),
.\key<129>.PAD.PAD (\key<129>.PAD.PAD ),
.\key<30>.PAD.PAD (\key<30>.PAD.PAD ),
.\key<179>.PAD.PAD (\key<179>.PAD.PAD ),
.\key<2>.PAD.PAD (\key<2>.PAD.PAD ),
.\key<50>.PAD.PAD (\key<50>.PAD.PAD ),
.\global_reset.PAD.PAD (\global_reset.PAD.PAD ),
.\key<64>.PAD.PAD (\key<64>.PAD.PAD ),
.\key<43>.PAD.PAD (\key<43>.PAD.PAD ),
.\key<214>.PAD.PAD (\key<214>.PAD.PAD ),
.\key<224>.PAD.PAD (\key<224>.PAD.PAD ),
.\encrypt<0>.PAD.PAD (\encrypt<0>.PAD.PAD ),
.\key<3>.PAD.PAD (\key<3>.PAD.PAD ),
.\key<63>.PAD.PAD (\key<63>.PAD.PAD ),
.\key<57>.PAD.PAD (\key<57>.PAD.PAD ),
.\count<0>.PAD.PAD (\count<0>.PAD.PAD ),
.\key<217>.PAD.PAD (\key<217>.PAD.PAD ),
.\key<66>.PAD.PAD (\key<66>.PAD.PAD ),
.\key<237>.PAD.PAD (\key<237>.PAD.PAD ),
.\key<56>.PAD.PAD (\key<56>.PAD.PAD ),
.\count<1>.PAD.PAD (\count<1>.PAD.PAD ),
.\key<216>.PAD.PAD (\key<216>.PAD.PAD ),
.\key<65>.PAD.PAD (\key<65>.PAD.PAD ),
.\key<236>.PAD.PAD (\key<236>.PAD.PAD ),
.\key<55>.PAD.PAD (\key<55>.PAD.PAD ),
.\key<229>.PAD.PAD (\key<229>.PAD.PAD ),
.\key<40>.PAD.PAD (\key<40>.PAD.PAD ),
.\key<69>.PAD.PAD (\key<69>.PAD.PAD ),
.\key<219>.PAD.PAD (\key<219>.PAD.PAD ),
.\key<239>.PAD.PAD (\key<239>.PAD.PAD ),
.\key<54>.PAD.PAD (\key<54>.PAD.PAD ),
.\key<249>.PAD.PAD (\key<249>.PAD.PAD ),
.\start<0>.PAD.PAD (\start<0>.PAD.PAD ),
.\my_clk.PAD.PAD (\my_clk.PAD.PAD ),
.\key<228>.PAD.PAD (\key<228>.PAD.PAD ),
.\key<68>.PAD.PAD (\key<68>.PAD.PAD ),
.\key<218>.PAD.PAD (\key<218>.PAD.PAD ),
.\key<238>.PAD.PAD (\key<238>.PAD.PAD ),
.\key<67>.PAD.PAD (\key<67>.PAD.PAD ),
.\key<248>.PAD.PAD (\key<248>.PAD.PAD ),
.\key<53>.PAD.PAD (\key<53>.PAD.PAD ),
.\key<208>.PAD.PAD (\key<208>.PAD.PAD ),
.\key<244>.PAD.PAD (\key<244>.PAD.PAD ),
.\key<132>.PAD.PAD (\key<132>.PAD.PAD ),
.\key<230>.PAD.PAD (\key<230>.PAD.PAD ),
.\key<146>.PAD.PAD (\key<146>.PAD.PAD ),
.\key<245>.PAD.PAD (\key<245>.PAD.PAD ),
.\key<209>.PAD.PAD (\key<209>.PAD.PAD ),
.\key<159>.PAD.PAD (\key<159>.PAD.PAD ),
.\key<131>.PAD.PAD (\key<131>.PAD.PAD ),
.\key<231>.PAD.PAD (\key<231>.PAD.PAD ),
.\key<145>.PAD.PAD (\key<145>.PAD.PAD ),
.\key<246>.PAD.PAD (\key<246>.PAD.PAD ),
.\key<134>.PAD.PAD (\key<134>.PAD.PAD ),
.\key<144>.PAD.PAD (\key<144>.PAD.PAD ),
.\key<247>.PAD.PAD (\key<247>.PAD.PAD ),
.\key<133>.PAD.PAD (\key<133>.PAD.PAD ),
.\key<143>.PAD.PAD (\key<143>.PAD.PAD ),
.\key<156>.PAD.PAD (\key<156>.PAD.PAD ),
.\key<254>.PAD.PAD (\key<254>.PAD.PAD ),
.\count<3>.PAD.PAD (\count<3>.PAD.PAD ),
.\key<240>.PAD.PAD (\key<240>.PAD.PAD ),
.\key<220>.PAD.PAD (\key<220>.PAD.PAD ),
.\key<136>.PAD.PAD (\key<136>.PAD.PAD ),
.\key<234>.PAD.PAD (\key<234>.PAD.PAD ),
.\key<155>.PAD.PAD (\key<155>.PAD.PAD ),
.\key<169>.PAD.PAD (\key<169>.PAD.PAD ),
.\key<255>.PAD.PAD (\key<255>.PAD.PAD ),
.\count<2>.PAD.PAD (\count<2>.PAD.PAD ),
.\key<241>.PAD.PAD (\key<241>.PAD.PAD ),
.\key<221>.PAD.PAD (\key<221>.PAD.PAD ),
.\key<235>.PAD.PAD (\key<235>.PAD.PAD ),
.\key<20>.PAD.PAD (\key<20>.PAD.PAD ),
.\key<149>.PAD.PAD (\key<149>.PAD.PAD ),
.\key<135>.PAD.PAD (\key<135>.PAD.PAD ),
.\key<252>.PAD.PAD (\key<252>.PAD.PAD ),
.\key<168>.PAD.PAD (\key<168>.PAD.PAD ),
.\key<158>.PAD.PAD (\key<158>.PAD.PAD ),
.\key<242>.PAD.PAD (\key<242>.PAD.PAD ),
.\key<138>.PAD.PAD (\key<138>.PAD.PAD ),
.\key<222>.PAD.PAD (\key<222>.PAD.PAD ),
.\key<232>.PAD.PAD (\key<232>.PAD.PAD ),
.\key<148>.PAD.PAD (\key<148>.PAD.PAD ),
.\key<253>.PAD.PAD (\key<253>.PAD.PAD ),
.\key<60>.PAD.PAD (\key<60>.PAD.PAD ),
.\key<157>.PAD.PAD (\key<157>.PAD.PAD ),
.\key<167>.PAD.PAD (\key<167>.PAD.PAD ),
.\key<243>.PAD.PAD (\key<243>.PAD.PAD ),
.\key<137>.PAD.PAD (\key<137>.PAD.PAD ),
.\key<223>.PAD.PAD (\key<223>.PAD.PAD ),
.\key<233>.PAD.PAD (\key<233>.PAD.PAD ),
.\key<147>.PAD.PAD (\key<147>.PAD.PAD ),
.\key<111>.PAD.PAD (\key<111>.PAD.PAD ),
.\key<125>.PAD.PAD (\key<125>.PAD.PAD ),
.\key<92>.PAD.PAD (\key<92>.PAD.PAD ),
.\key<194>.PAD.PAD (\key<194>.PAD.PAD ),
.\key<23>.PAD.PAD (\key<23>.PAD.PAD ),
.\key<24>.PAD.PAD (\key<24>.PAD.PAD ),
.\key<82>.PAD.PAD (\key<82>.PAD.PAD ),
.\key<166>.PAD.PAD (\key<166>.PAD.PAD ),
.\key<250>.PAD.PAD (\key<250>.PAD.PAD ),
.\key<200>.PAD.PAD (\key<200>.PAD.PAD ),
.\key<72>.PAD.PAD (\key<72>.PAD.PAD ),
.\key<152>.PAD.PAD (\key<152>.PAD.PAD ),
.\key<10>.PAD.PAD (\key<10>.PAD.PAD ),
.\key<112>.PAD.PAD (\key<112>.PAD.PAD ),
.\key<91>.PAD.PAD (\key<91>.PAD.PAD ),
.\key<126>.PAD.PAD (\key<126>.PAD.PAD ),
.\key<193>.PAD.PAD (\key<193>.PAD.PAD ),
.\key<25>.PAD.PAD (\key<25>.PAD.PAD ),
.\key<165>.PAD.PAD (\key<165>.PAD.PAD ),
.\key<201>.PAD.PAD (\key<201>.PAD.PAD ),
.\key<251>.PAD.PAD (\key<251>.PAD.PAD ),
.\key<81>.PAD.PAD (\key<81>.PAD.PAD ),
.\key<71>.PAD.PAD (\key<71>.PAD.PAD ),
.\key<151>.PAD.PAD (\key<151>.PAD.PAD ),
.\key<123>.PAD.PAD (\key<123>.PAD.PAD ),
.\key<11>.PAD.PAD (\key<11>.PAD.PAD ),
.\key<21>.PAD.PAD (\key<21>.PAD.PAD ),
.\key<90>.PAD.PAD (\key<90>.PAD.PAD ),
.\key<113>.PAD.PAD (\key<113>.PAD.PAD ),
.\key<202>.PAD.PAD (\key<202>.PAD.PAD ),
.\key<192>.PAD.PAD (\key<192>.PAD.PAD ),
.\key<84>.PAD.PAD (\key<84>.PAD.PAD ),
.\key<164>.PAD.PAD (\key<164>.PAD.PAD ),
.\key<70>.PAD.PAD (\key<70>.PAD.PAD ),
.\key<154>.PAD.PAD (\key<154>.PAD.PAD ),
.\key<124>.PAD.PAD (\key<124>.PAD.PAD ),
.\key<114>.PAD.PAD (\key<114>.PAD.PAD ),
.\key<12>.PAD.PAD (\key<12>.PAD.PAD ),
.\key<22>.PAD.PAD (\key<22>.PAD.PAD ),
.\key<203>.PAD.PAD (\key<203>.PAD.PAD ),
.\key<163>.PAD.PAD (\key<163>.PAD.PAD ),
.\key<191>.PAD.PAD (\key<191>.PAD.PAD ),
.\key<83>.PAD.PAD (\key<83>.PAD.PAD ),
.\key<153>.PAD.PAD (\key<153>.PAD.PAD ),
.\key<13>.PAD.PAD (\key<13>.PAD.PAD ),
.\key<170>.PAD.PAD (\key<170>.PAD.PAD ),
.\key<142>.PAD.PAD (\key<142>.PAD.PAD ),
.\key<121>.PAD.PAD (\key<121>.PAD.PAD ),
.\key<180>.PAD.PAD (\key<180>.PAD.PAD ),
.\key<96>.PAD.PAD (\key<96>.PAD.PAD ),
.\key<14>.PAD.PAD (\key<14>.PAD.PAD ),
.\key<101>.PAD.PAD (\key<101>.PAD.PAD ),
.\key<162>.PAD.PAD (\key<162>.PAD.PAD ),
.\key<190>.PAD.PAD (\key<190>.PAD.PAD ),
.\key<28>.PAD.PAD (\key<28>.PAD.PAD ),
.\key<204>.PAD.PAD (\key<204>.PAD.PAD ),
.\key<141>.PAD.PAD (\key<141>.PAD.PAD ),
.\key<95>.PAD.PAD (\key<95>.PAD.PAD ),
.\key<122>.PAD.PAD (\key<122>.PAD.PAD ),
.\key<102>.PAD.PAD (\key<102>.PAD.PAD ),
.\key<15>.PAD.PAD (\key<15>.PAD.PAD ),
.\key<161>.PAD.PAD (\key<161>.PAD.PAD ),
.\key<205>.PAD.PAD (\key<205>.PAD.PAD ),
.\key<29>.PAD.PAD (\key<29>.PAD.PAD ),
.\key<160>.PAD.PAD (\key<160>.PAD.PAD ),
.\key<140>.PAD.PAD (\key<140>.PAD.PAD ),
.\key<94>.PAD.PAD (\key<94>.PAD.PAD ),
.\key<130>.PAD.PAD (\key<130>.PAD.PAD ),
.\key<182>.PAD.PAD (\key<182>.PAD.PAD ),
.\key<150>.PAD.PAD (\key<150>.PAD.PAD ),
.\key<16>.PAD.PAD (\key<16>.PAD.PAD ),
.\key<80>.PAD.PAD (\key<80>.PAD.PAD ),
.\key<206>.PAD.PAD (\key<206>.PAD.PAD ),
.\key<26>.PAD.PAD (\key<26>.PAD.PAD ),
.\key<110>.PAD.PAD (\key<110>.PAD.PAD ),
.\key<181>.PAD.PAD (\key<181>.PAD.PAD ),
.\key<93>.PAD.PAD (\key<93>.PAD.PAD ),
.\key<120>.PAD.PAD (\key<120>.PAD.PAD ),
.\key<100>.PAD.PAD (\key<100>.PAD.PAD ),
.\key<17>.PAD.PAD (\key<17>.PAD.PAD ),
.\key<27>.PAD.PAD (\key<27>.PAD.PAD ),
.\key<207>.PAD.PAD (\key<207>.PAD.PAD ),
.\KSi<19>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<19>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<163>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<163>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<17>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<17>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<55>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<55>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<37>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<37>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<26>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<26>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<136>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<136>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<174>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<174>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<67>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<67>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<6>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<6>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<77>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<77>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<15>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<15>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<108>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<108>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<13>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<13>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<86>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<86>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<150>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<150>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<85>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<85>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<157>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<157>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<113>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<113>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<41>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<41>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<110>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<110>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<104>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<104>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<83>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<83>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<89>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<89>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<11>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<11>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<7>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<7>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<164>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<164>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<179>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<179>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<109>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<109>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<173>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<173>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<155>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<155>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<31>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<31>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<123>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<123>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<44>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<44>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<84>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<84>_FINAL_OUTPUT.OUTBUF.OUT ),
.\new_count<2>_FINAL_OUTPUT.OUTBUF.OUT (\new_count<2>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<5>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<5>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<118>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<118>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<141>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<141>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<165>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<165>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<130>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<130>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<162>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<162>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<33>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<33>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<161>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<161>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<154>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<154>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<64>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<64>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<78>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<78>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<170>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<170>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<1>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<1>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<135>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<135>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<95>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<95>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<139>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<139>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<49>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<49>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<12>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<12>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<146>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<146>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<61>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<61>_FINAL_OUTPUT.OUTBUF.OUT ),
.\data_ready<0>_FINAL_OUTPUT.OUTBUF.OUT (\data_ready<0>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<34>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<34>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<62>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<62>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<24>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<24>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<53>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<53>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<0>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<0>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<125>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<125>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<22>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<22>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<9>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<9>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<48>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<48>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<111>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<111>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<70>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<70>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<74>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<74>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<79>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<79>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<58>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<58>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<2>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<2>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<29>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<29>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<148>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<148>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<186>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<186>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<68>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<68>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<99>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<99>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<190>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<190>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<105>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<105>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<119>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<119>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<35>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<35>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<133>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<133>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<188>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<188>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<158>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<158>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<115>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<115>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<46>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<46>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<93>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<93>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<73>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<73>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<28>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<28>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<143>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<143>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<54>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<54>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<18>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<18>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<177>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<177>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<106>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<106>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<98>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<98>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<30>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<30>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<142>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<142>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<167>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<167>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<3>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<3>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<60>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<60>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<181>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<181>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<39>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<39>_FINAL_OUTPUT.OUTBUF.OUT ),
.\new_count<0>_FINAL_OUTPUT.OUTBUF.OUT (\new_count<0>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<132>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<132>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<16>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<16>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<191>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<191>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<45>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<45>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<116>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<116>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<47>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<47>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<81>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<81>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<100>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<100>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<168>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<168>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<59>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<59>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<121>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<121>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<72>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<72>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<159>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<159>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<14>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<14>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<25>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<25>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<82>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<82>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<90>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<90>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<36>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<36>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<97>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<97>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<175>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<175>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<134>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<134>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<151>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<151>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<10>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<10>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<80>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<80>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<138>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<138>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<169>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<169>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<149>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<149>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<176>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<176>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<140>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<140>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<71>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<71>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<153>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<153>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<145>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<145>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<124>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<124>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<8>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<8>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<172>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<172>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<40>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<40>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<96>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<96>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<75>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<75>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<103>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<103>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<122>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<122>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<129>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<129>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<183>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<183>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<156>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<156>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<4>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<4>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<38>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<38>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<128>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<128>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<107>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<107>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<23>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<23>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<88>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<88>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<185>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<185>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<57>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<57>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<187>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<187>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<50>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<50>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<160>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<160>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<144>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<144>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<32>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<32>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<21>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<21>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<102>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<102>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<137>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<137>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<131>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<131>_FINAL_OUTPUT.OUTBUF.OUT ),
.\new_count<1>_FINAL_OUTPUT.OUTBUF.OUT (\new_count<1>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<152>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<152>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<94>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<94>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<182>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<182>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<189>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<189>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<56>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<56>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<52>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<52>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<171>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<171>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<87>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<87>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<51>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<51>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<65>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<65>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<114>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<114>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<76>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<76>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<126>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<126>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<91>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<91>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<92>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<92>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<117>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<117>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<27>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<27>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<66>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<66>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<69>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<69>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<101>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<101>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<178>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<178>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<43>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<43>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<112>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<112>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<166>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<166>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<180>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<180>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<127>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<127>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<147>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<147>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<184>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<184>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<20>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<20>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<42>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<42>_FINAL_OUTPUT.OUTBUF.OUT ),
.\new_count<3>_FINAL_OUTPUT.OUTBUF.OUT (\new_count<3>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<120>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<120>_FINAL_OUTPUT.OUTBUF.OUT ),
.\KSi<63>_FINAL_OUTPUT.OUTBUF.OUT (\KSi<63>_FINAL_OUTPUT.OUTBUF.OUT )
);

initial begin
// Initialize Inputs
\key<173>.PAD.PAD  = 0;
\key<89>.PAD.PAD  = 0;
\key<8>.PAD.PAD  = 0;
\key<183>.PAD.PAD  = 0;
\key<108>.PAD.PAD  = 0;
\key<99>.PAD.PAD  = 0;
\key<174>.PAD.PAD  = 0;
\key<9>.PAD.PAD  = 0;
\key<184>.PAD.PAD  = 0;
\key<107>.PAD.PAD  = 0;
\key<39>.PAD.PAD  = 0;
\key<19>.PAD.PAD  = 0;
\key<77>.PAD.PAD  = 0;
\key<185>.PAD.PAD  = 0;
\key<97>.PAD.PAD  = 0;
\key<199>.PAD.PAD  = 0;
\key<171>.PAD.PAD  = 0;
\key<59>.PAD.PAD  = 0;
\key<38>.PAD.PAD  = 0;
\key<172>.PAD.PAD  = 0;
\key<18>.PAD.PAD  = 0;
\key<78>.PAD.PAD  = 0;
\key<186>.PAD.PAD  = 0;
\key<109>.PAD.PAD  = 0;
\key<98>.PAD.PAD  = 0;
\key<79>.PAD.PAD  = 0;
\key<119>.PAD.PAD  = 0;
\key<58>.PAD.PAD  = 0;
\key<187>.PAD.PAD  = 0;
\key<47>.PAD.PAD  = 0;
\key<75>.PAD.PAD  = 0;
\key<4>.PAD.PAD  = 0;
\key<37>.PAD.PAD  = 0;
\key<177>.PAD.PAD  = 0;
\key<85>.PAD.PAD  = 0;
\key<118>.PAD.PAD  = 0;
\key<197>.PAD.PAD  = 0;
\key<104>.PAD.PAD  = 0;
\key<188>.PAD.PAD  = 0;
\key<5>.PAD.PAD  = 0;
\key<76>.PAD.PAD  = 0;
\key<46>.PAD.PAD  = 0;
\key<36>.PAD.PAD  = 0;
\key<86>.PAD.PAD  = 0;
\key<178>.PAD.PAD  = 0;
\key<117>.PAD.PAD  = 0;
\key<198>.PAD.PAD  = 0;
\key<45>.PAD.PAD  = 0;
\key<103>.PAD.PAD  = 0;
\key<6>.PAD.PAD  = 0;
\key<49>.PAD.PAD  = 0;
\key<211>.PAD.PAD  = 0;
\key<73>.PAD.PAD  = 0;
\key<189>.PAD.PAD  = 0;
\key<87>.PAD.PAD  = 0;
\key<35>.PAD.PAD  = 0;
\key<175>.PAD.PAD  = 0;
\key<116>.PAD.PAD  = 0;
\key<34>.PAD.PAD  = 0;
\key<195>.PAD.PAD  = 0;
\key<106>.PAD.PAD  = 0;
\key<48>.PAD.PAD  = 0;
\key<7>.PAD.PAD  = 0;
\key<210>.PAD.PAD  = 0;
\key<74>.PAD.PAD  = 0;
\key<176>.PAD.PAD  = 0;
\key<88>.PAD.PAD  = 0;
\key<33>.PAD.PAD  = 0;
\key<115>.PAD.PAD  = 0;
\key<196>.PAD.PAD  = 0;
\key<105>.PAD.PAD  = 0;
\key<213>.PAD.PAD  = 0;
\key<42>.PAD.PAD  = 0;
\key<127>.PAD.PAD  = 0;
\key<32>.PAD.PAD  = 0;
\key<227>.PAD.PAD  = 0;
\key<0>.PAD.PAD  = 0;
\key<52>.PAD.PAD  = 0;
\key<62>.PAD.PAD  = 0;
\key<41>.PAD.PAD  = 0;
\key<128>.PAD.PAD  = 0;
\key<226>.PAD.PAD  = 0;
\key<31>.PAD.PAD  = 0;
\key<212>.PAD.PAD  = 0;
\key<1>.PAD.PAD  = 0;
\key<51>.PAD.PAD  = 0;
\key<61>.PAD.PAD  = 0;
\key<139>.PAD.PAD  = 0;
\key<44>.PAD.PAD  = 0;
\key<215>.PAD.PAD  = 0;
\key<225>.PAD.PAD  = 0;
\key<129>.PAD.PAD  = 0;
\key<30>.PAD.PAD  = 0;
\key<179>.PAD.PAD  = 0;
\key<2>.PAD.PAD  = 0;
\key<50>.PAD.PAD  = 0;
\global_reset.PAD.PAD  = 0;
\key<64>.PAD.PAD  = 0;
\key<43>.PAD.PAD  = 0;
\key<214>.PAD.PAD  = 0;
\key<224>.PAD.PAD  = 0;
\encrypt<0>.PAD.PAD  = 0;
\key<3>.PAD.PAD  = 0;
\key<63>.PAD.PAD  = 0;
\key<57>.PAD.PAD  = 0;
\count<0>.PAD.PAD  = 0;
\key<217>.PAD.PAD  = 0;
\key<66>.PAD.PAD  = 0;
\key<237>.PAD.PAD  = 0;
\key<56>.PAD.PAD  = 0;
\count<1>.PAD.PAD  = 0;
\key<216>.PAD.PAD  = 0;
\key<65>.PAD.PAD  = 0;
\key<236>.PAD.PAD  = 0;
\key<55>.PAD.PAD  = 0;
\key<229>.PAD.PAD  = 0;
\key<40>.PAD.PAD  = 0;
\key<69>.PAD.PAD  = 0;
\key<219>.PAD.PAD  = 0;
\key<239>.PAD.PAD  = 0;
\key<54>.PAD.PAD  = 0;
\key<249>.PAD.PAD  = 0;
\start<0>.PAD.PAD  = 0;
\my_clk.PAD.PAD  = 0;
\key<228>.PAD.PAD  = 0;
\key<68>.PAD.PAD  = 0;
\key<218>.PAD.PAD  = 0;
\key<238>.PAD.PAD  = 0;
\key<67>.PAD.PAD  = 0;
\key<248>.PAD.PAD  = 0;
\key<53>.PAD.PAD  = 0;
\key<208>.PAD.PAD  = 0;
\key<244>.PAD.PAD  = 0;
\key<132>.PAD.PAD  = 0;
\key<230>.PAD.PAD  = 0;
\key<146>.PAD.PAD  = 0;
\key<245>.PAD.PAD  = 0;
\key<209>.PAD.PAD  = 0;
\key<159>.PAD.PAD  = 0;
\key<131>.PAD.PAD  = 0;
\key<231>.PAD.PAD  = 0;
\key<145>.PAD.PAD  = 0;
\key<246>.PAD.PAD  = 0;
\key<134>.PAD.PAD  = 0;
\key<144>.PAD.PAD  = 0;
\key<247>.PAD.PAD  = 0;
\key<133>.PAD.PAD  = 0;
\key<143>.PAD.PAD  = 0;
\key<156>.PAD.PAD  = 0;
\key<254>.PAD.PAD  = 0;
\count<3>.PAD.PAD  = 0;
\key<240>.PAD.PAD  = 0;
\key<220>.PAD.PAD  = 0;
\key<136>.PAD.PAD  = 0;
\key<234>.PAD.PAD  = 0;
\key<155>.PAD.PAD  = 0;
\key<169>.PAD.PAD  = 0;
\key<255>.PAD.PAD  = 0;
\count<2>.PAD.PAD  = 0;
\key<241>.PAD.PAD  = 0;
\key<221>.PAD.PAD  = 0;
\key<235>.PAD.PAD  = 0;
\key<20>.PAD.PAD  = 0;
\key<149>.PAD.PAD  = 0;
\key<135>.PAD.PAD  = 0;
\key<252>.PAD.PAD  = 0;
\key<168>.PAD.PAD  = 0;
\key<158>.PAD.PAD  = 0;
\key<242>.PAD.PAD  = 0;
\key<138>.PAD.PAD  = 0;
\key<222>.PAD.PAD  = 0;
\key<232>.PAD.PAD  = 0;
\key<148>.PAD.PAD  = 0;
\key<253>.PAD.PAD  = 0;
\key<60>.PAD.PAD  = 0;
\key<157>.PAD.PAD  = 0;
\key<167>.PAD.PAD  = 0;
\key<243>.PAD.PAD  = 0;
\key<137>.PAD.PAD  = 0;
\key<223>.PAD.PAD  = 0;
\key<233>.PAD.PAD  = 0;
\key<147>.PAD.PAD  = 0;
\key<111>.PAD.PAD  = 0;
\key<125>.PAD.PAD  = 0;
\key<92>.PAD.PAD  = 0;
\key<194>.PAD.PAD  = 0;
\key<23>.PAD.PAD  = 0;
\key<24>.PAD.PAD  = 0;
\key<82>.PAD.PAD  = 0;
\key<166>.PAD.PAD  = 0;
\key<250>.PAD.PAD  = 0;
\key<200>.PAD.PAD  = 0;
\key<72>.PAD.PAD  = 0;
\key<152>.PAD.PAD  = 0;
\key<10>.PAD.PAD  = 0;
\key<112>.PAD.PAD  = 0;
\key<91>.PAD.PAD  = 0;
\key<126>.PAD.PAD  = 0;
\key<193>.PAD.PAD  = 0;
\key<25>.PAD.PAD  = 0;
\key<165>.PAD.PAD  = 0;
\key<201>.PAD.PAD  = 0;
\key<251>.PAD.PAD  = 0;
\key<81>.PAD.PAD  = 0;
\key<71>.PAD.PAD  = 0;
\key<151>.PAD.PAD  = 0;
\key<123>.PAD.PAD  = 0;
\key<11>.PAD.PAD  = 0;
\key<21>.PAD.PAD  = 0;
\key<90>.PAD.PAD  = 0;
\key<113>.PAD.PAD  = 0;
\key<202>.PAD.PAD  = 0;
\key<192>.PAD.PAD  = 0;
\key<84>.PAD.PAD  = 0;
\key<164>.PAD.PAD  = 0;
\key<70>.PAD.PAD  = 0;
\key<154>.PAD.PAD  = 0;
\key<124>.PAD.PAD  = 0;
\key<114>.PAD.PAD  = 0;
\key<12>.PAD.PAD  = 0;
\key<22>.PAD.PAD  = 0;
\key<203>.PAD.PAD  = 0;
\key<163>.PAD.PAD  = 0;
\key<191>.PAD.PAD  = 0;
\key<83>.PAD.PAD  = 0;
\key<153>.PAD.PAD  = 0;
\key<13>.PAD.PAD  = 0;
\key<170>.PAD.PAD  = 0;
\key<142>.PAD.PAD  = 0;
\key<121>.PAD.PAD  = 0;
\key<180>.PAD.PAD  = 0;
\key<96>.PAD.PAD  = 0;
\key<14>.PAD.PAD  = 0;
\key<101>.PAD.PAD  = 0;
\key<162>.PAD.PAD  = 0;
\key<190>.PAD.PAD  = 0;
\key<28>.PAD.PAD  = 0;
\key<204>.PAD.PAD  = 0;
\key<141>.PAD.PAD  = 0;
\key<95>.PAD.PAD  = 0;
\key<122>.PAD.PAD  = 0;
\key<102>.PAD.PAD  = 0;
\key<15>.PAD.PAD  = 0;
\key<161>.PAD.PAD  = 0;
\key<205>.PAD.PAD  = 0;
\key<29>.PAD.PAD  = 0;
\key<160>.PAD.PAD  = 0;
\key<140>.PAD.PAD  = 0;
\key<94>.PAD.PAD  = 0;
\key<130>.PAD.PAD  = 0;
\key<182>.PAD.PAD  = 0;
\key<150>.PAD.PAD  = 0;
\key<16>.PAD.PAD  = 0;
\key<80>.PAD.PAD  = 0;
\key<206>.PAD.PAD  = 0;
\key<26>.PAD.PAD  = 0;
\key<110>.PAD.PAD  = 0;
\key<181>.PAD.PAD  = 0;
\key<93>.PAD.PAD  = 0;
\key<120>.PAD.PAD  = 0;
\key<100>.PAD.PAD  = 0;
\key<17>.PAD.PAD  = 0;
\key<27>.PAD.PAD  = 0;
\key<207>.PAD.PAD  = 0;


// Wait 100 ns for global reset to finish
	#100;

	// Add stimulus here

end

endmodule