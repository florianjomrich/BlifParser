`timescale 1ns / 1ps 
 
module TEST; 
 
// Inputs 
reg \in1.PAD.PAD ;
reg \newCLK.PAD.PAD ;
reg \global_reset.PAD.PAD ;

// Outputs 
wire \out6_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out9_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out11_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out14_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out8_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out15_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out7_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out1_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out13_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out12_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out5_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out10_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out2_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out3_FINAL_OUTPUT.OUTBUF.OUT ;
wire \out4_FINAL_OUTPUT.OUTBUF.OUT ;
 
// Instantiate the Unit Under Test (UUT) 
 
HelloWorld uut (
.\in1.PAD.PAD (\in1.PAD.PAD ),
.\newCLK.PAD.PAD (\newCLK.PAD.PAD ),
.\global_reset.PAD.PAD (\global_reset.PAD.PAD ),
.\out6_FINAL_OUTPUT.OUTBUF.OUT (\out6_FINAL_OUTPUT.OUTBUF.OUT ),
.\out9_FINAL_OUTPUT.OUTBUF.OUT (\out9_FINAL_OUTPUT.OUTBUF.OUT ),
.\out11_FINAL_OUTPUT.OUTBUF.OUT (\out11_FINAL_OUTPUT.OUTBUF.OUT ),
.\out14_FINAL_OUTPUT.OUTBUF.OUT (\out14_FINAL_OUTPUT.OUTBUF.OUT ),
.\out8_FINAL_OUTPUT.OUTBUF.OUT (\out8_FINAL_OUTPUT.OUTBUF.OUT ),
.\out15_FINAL_OUTPUT.OUTBUF.OUT (\out15_FINAL_OUTPUT.OUTBUF.OUT ),
.\out7_FINAL_OUTPUT.OUTBUF.OUT (\out7_FINAL_OUTPUT.OUTBUF.OUT ),
.\out1_FINAL_OUTPUT.OUTBUF.OUT (\out1_FINAL_OUTPUT.OUTBUF.OUT ),
.\out13_FINAL_OUTPUT.OUTBUF.OUT (\out13_FINAL_OUTPUT.OUTBUF.OUT ),
.\out12_FINAL_OUTPUT.OUTBUF.OUT (\out12_FINAL_OUTPUT.OUTBUF.OUT ),
.\out5_FINAL_OUTPUT.OUTBUF.OUT (\out5_FINAL_OUTPUT.OUTBUF.OUT ),
.\out10_FINAL_OUTPUT.OUTBUF.OUT (\out10_FINAL_OUTPUT.OUTBUF.OUT ),
.\out2_FINAL_OUTPUT.OUTBUF.OUT (\out2_FINAL_OUTPUT.OUTBUF.OUT ),
.\out3_FINAL_OUTPUT.OUTBUF.OUT (\out3_FINAL_OUTPUT.OUTBUF.OUT ),
.\out4_FINAL_OUTPUT.OUTBUF.OUT (\out4_FINAL_OUTPUT.OUTBUF.OUT )
);

initial begin
// Initialize Inputs
\in1.PAD.PAD  = 0;
\newCLK.PAD.PAD  = 0;
\global_reset.PAD.PAD  = 0;


// Wait 100 ns for global reset to finish
	#100;

	// Add stimulus here

end

endmodule