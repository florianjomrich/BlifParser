//    Xilinx Proprietary Primitive Cell X_ZERO for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verplex_libs/data/simprims/X_ZERO.v,v 1.4.198.3 2004/09/28 20:47:47 wloo Exp $
//

`celldefine
`timescale 1 ps/1 ps

module X_ZERO (O);

  output O;

  assign O = 1'b0;

endmodule
