//    Xilinx Proprietary Primitive Cell X_SUH for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verplex_libs/data/simprims/X_SUH.v,v 1.3.198.3 2004/09/28 20:47:46 wloo Exp $
//

`celldefine
`timescale 1 ps/1 ps

module X_SUH (I, CE, CLK);

  input I, CLK, CE;

endmodule
