//    Xilinx Proprietary Primitive Cell X_BPAD for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verplex_libs/data/simprims/X_BPAD.v,v 1.3.198.3 2004/09/28 20:47:45 wloo Exp $
//

`celldefine
`timescale 1 ps/1 ps

module X_BPAD (PAD);

  input PAD;

endmodule
