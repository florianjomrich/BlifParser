// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verplex_libs/data/simprims/Attic/X_IDELAYCTRL.v,v 1.1.2.1 2004/09/28 20:47:46 wloo Exp $

`timescale 1 ps / 1 ps 

module X_IDELAYCTRL (RDY, REFCLK, RST);

    output RDY;
    input REFCLK;
    input RST;

endmodule // X_IDELAYCTRL
